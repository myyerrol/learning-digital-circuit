module mst_3(
);

endmodule
